---------------------------------------------------------------------------------
--
-- Copyright (c) 2017 by SISLAB Team, LSI Design Contest 2018.
-- The University of Engineering and Technology, Vietnam National University.
-- All right resevered.
--
-- Copyright notification
-- No part may be reproduced except as authorized by written permission.
-- 
-- @File            : !!FILE
-- @Author          : Van-Nam DINH       @Modifier      : Van-Nam DINH
-- @Created Date    : !!DATE       @Modified Date : !!DATE
-- @Project         : Artificial Neural Network
-- @Module          : !!MODULE
-- @Description     :
-- @Version         :
-- @ID              :
--
---------------------------------------------------------------------------------

---------------------------------------------------------------------------------
-- Library declaration
---------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

---------------------------------------------------------------------------------
-- Entity declaration
--------------------------------------------------------------------------------- 
entity !!MODULE is
    port(
        clk     : in std_logic;
        rst     : in std_logic;
    );
end entity; 

---------------------------------------------------------------------------------
-- Architecture description
---------------------------------------------------------------------------------
architecture behavior of !!MODULE is
  
begin

end behavior;
