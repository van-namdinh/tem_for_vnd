--------------------------------------------------------------------------------
-- Project name   :
-- File name      : !!FILE
-- Created date   : !!DATE
-- Author         : Huy-Hung Ho
-- Last modified  : !!DATE
-- Desc           :
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity  is
    port {
    
    }
end entity;

architecture behavior of  is

begin

end;
